//`include "CoreTest.sv"
`include "ControllerTest.sv"
