//`include "core_test.sv"
`include "controllerTest.sv"
//`include "types_test.sv"
