`include "core_test.sv"
//`include "types_test.sv"
