`include "BusInterface.svh"

module Controller #(
  parameter 	p_WIDTH = 32
) (
  BusInterface.controller intf
);

endmodule